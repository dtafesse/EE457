LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;


entity de1_top is
generic (
  simulation_wide : positive := 28;    -- used for simulation to overide width
  simulation_max  : positive := 50000000); -- used for simulaiton to oreride max value
port
(
	-- 50Mhz clock, i.e. 50 Million rising edges per second
   clock_50 :in  std_logic; 
    -- 7 Segment Display
	hex0     :out std_logic_vector(6 downto 0); -- right most
	hex1     :out std_logic_vector(6 downto 0);	
	hex2     :out std_logic_vector(6 downto 0);	
	hex3     :out std_logic_vector(6 downto 0);	
	hex4     :out std_logic_vector(6 downto 0);	
	hex5     :out std_logic_vector(6 downto 0); -- left most
    -- Red LEDs above Slider switches
	-- drive the ledr's high to light them up
    ledr     :out std_logic_vector(9 downto 0);
	-- key/Push Button, push button to drive a signal low, normally high
	key      :in  std_logic_vector(3 downto 0);  
    -- Slider Switch, logic 0 when slide down, logic 1 when pushed towards 7 segments
	sw       :in	 std_logic_vector(9 downto 0) 
);

end de1_top;

architecture struct of de1_top is

-- define signals to be used
signal enable_pulse_every_second     : std_logic;
signal reset_n                       : std_logic;
signal one_second_count_value        : std_logic_vector(3 downto 0);
signal ten_second_count_value        : std_logic_vector(3 downto 0);
signal enable_pulse_every_10_second  : std_logic;
signal load_counter                  : std_logic;


-- define the component
component gen_counter is
generic (
		wide :positive; -- how many bits is the counter
		max  :positive  -- what is the max count
		);
port (
		clk	     :in	std_logic;
		data	 :in  std_logic_vector(wide-1 downto 0 );
		load	 :in  std_logic;
		enable   :in  std_logic;
		reset_n	 :in  std_logic;
		count	 :out std_logic_vector(wide-1 downto 0 );
		term	 :out std_logic);
	end component;
	

component seven_segment_cntrl IS
	-- Begin port declaration
	port (
		-- Declare data input "input"
		input : in unsigned(3 downto 0);
		-- Declare the seven segment output
		hex   : out std_logic_vector(6 downto 0));
-- End entity		
end component;

begin

-- turn off the other 7 segments, drive high to turn off
--hex1 <= (others => '1');
hex2 <= (others => '1');
hex3 <= (others => '1');
hex4 <= (others => '1');
hex5 <= (others => '1');

-- turn off unused LEDs, drive 0 to keep off
--ledr(7 downto 4) <= (others =>'0');


-- use a name that makes sense, key(0) is our reset, push to reset
reset_n <= key(0);  -- key is normally high


-- first use an instance of counter to get clock enable
-- never ever use the term output as clock, always use as an enable 
large_counter : gen_counter
generic map (
		wide => simulation_wide, -- need 28 bits do divide 50Mhz down to 1 second
		max  => simulation_max   -- terminate the count when you hit 50Million
		)
port map (
		clk      => clock_50,
		data	 => (others => '0'),
		load	 => '0',   -- not loadable
		enable   => '1',   -- always enabled
		reset_n	 => reset_n, 
		count	 => open,  -- we are not using this signal
		term	 => enable_pulse_every_second -- goes high for 1 clock cycle max value hit
		);
	
load_counter <= not key(1); -- need to invert, key is normally high		
-- this counter will count seconds.			
one_second_counter : gen_counter 
generic map (
		wide => 4,  -- created a 4 bit counter (max count could be 15)
		max  => 9   -- stop counting after 9, go back to 0
		)
port map (
		clk	     => clock_50,
		data	 => sw(3 downto 0), -- use switch for data input to preload
		load	 => load_counter,   
		enable   => enable_pulse_every_second,
		reset_n	 => reset_n,
		count	 => one_second_count_value,
		term	 => enable_pulse_every_10_second);-- this signal will pulse for 1 clock cycle when the cunter roles over
		
		
-- turn the LED 8 on when the terminal count has been hit, should be after 10 seconds
ledr(8) <=  enable_pulse_every_10_second;  
-- turn the LED 9 on when the terminal count for 1 second is hit, every 1 second
ledr(9) <=  enable_pulse_every_second;
-- question, why can't you see the above LEDs light up?

-- drive the value out the low 4 red leds
ledr(3 downto 0) <= one_second_count_value;
ledr(7 downto 4) <= ten_second_count_value;

ten_second_counter : gen_counter 
generic map (
		wide => 4,  -- created a 4 bit counter (max count would be 15)
		max  => 5   -- stop counting after 5, go back to 0
		)
port map (
		clk	     => clock_50,
		data	 => sw(7 downto 4), -- use switch for data input to preload
		load	 => load_counter,   
		enable   => enable_pulse_every_10_second,
		reset_n	 => reset_n,
		count	 => ten_second_count_value,
		term	 => open);


hex0_driver: seven_segment_cntrl
	-- Begin port declaration
  port map(
    input => unsigned(one_second_count_value),
	hex   => hex0); 

hex1_driver: seven_segment_cntrl
	-- Begin port declaration
  port map(
    input => unsigned(ten_second_count_value),
	hex   => hex1); 
	 
end; -- end the design









